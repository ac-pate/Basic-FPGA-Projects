library IEEE;
use IEEE.std_logic_1164.all;

entity sum_of_minterms is
port( a,b,c       : in std_logic;
output            : out std_logic);
end sum_of_minterms;
